`timescale 1ns / 1ps

module Core(
  input clk,
  input rst,
);

  //

endmodule // Core
